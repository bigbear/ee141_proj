** Generated for: hspiceD
** Generated on: Sep 17 17:04:59 2012
** Design library name: labs
** Design cell name: inv
** Design view name: extracted


.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    MEASOUT=1
+    PARHIER=LOCAL
+    PSF=2

** Library name: labs
** Cell name: inv
** View name: extracted
m0 out in vdd! vdd! gpdk090_pmos1v L=100e-9 W=240e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
m1 out in 0 0 gpdk090_nmos1v L=100e-9 W=120e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
.END
