** Generated for: hspiceD
** Generated on: Sep 24 14:59:14 2012
** Design library name: labs
** Design cell name: 5-stage_inv
** Design view name: extracted


.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    MEASOUT=1
+    PARHIER=LOCAL
+    PSF=2

** Library name: labs
** Cell name: 5-stage_inv
** View name: extracted
m0 n1 n5 n7 n7 gpdk090_pmos1v L=100e-9 W=240e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
m1 n5 n4 n7 n7 gpdk090_pmos1v L=100e-9 W=240e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
m2 n4 n3 n7 n7 gpdk090_pmos1v L=100e-9 W=240e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
m3 n3 n2 n7 n7 gpdk090_pmos1v L=100e-9 W=240e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
m4 n2 n1 n7 n7 gpdk090_pmos1v L=100e-9 W=240e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
m5 n1 n5 n6 n6 gpdk090_nmos1v L=100e-9 W=120e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
m6 n5 n4 n6 n6 gpdk090_nmos1v L=100e-9 W=120e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
m7 n4 n3 n6 n6 gpdk090_nmos1v L=100e-9 W=120e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
m8 n3 n2 n6 n6 gpdk090_nmos1v L=100e-9 W=120e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
m9 n2 n1 n6 n6 gpdk090_nmos1v L=100e-9 W=120e-9 AD=69.6e-15 AS=69.6e-15 PD=1.16e-6 PS=1.16e-6 M=1
.END
